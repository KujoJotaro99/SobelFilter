`timescale 1ns/1ps

module conv2d 
#(
    parameter WIDTH_P = 8,
    parameter DEPTH_P = 16
)(
    input  logic clk_i,
    input  logic rstn_i,
    input  logic valid_i,
    input  logic ready_i,
    input  logic [WIDTH_P-1:0] data_i,
    output logic valid_o,
    output logic ready_o,
    output logic signed [(2*WIDTH_P)-1:0] gx_o,
    output logic signed [(2*WIDTH_P)-1:0] gy_o
);

    logic [WIDTH_P-1:0] ram_row0, ram_row1;

    // likely need some kind of delayed valid with the ram because contents not cleared between test, only conv window is cleared so the circular buffer may dump wrong values
    ramdelaybuffer #(
        .WIDTH_P(WIDTH_P),
        .DELAY_P(2*DEPTH_P-1),
        .DELAY_A_P(2*DEPTH_P-1),
        .DELAY_B_P(DEPTH_P-1)
    ) line_buffer (
        .clk_i(clk_i),
        .rstn_i(rstn_i),
        .valid_i(valid_i),
        .ready_i(ready_i),
        .valid_o(valid_o),
        .ready_o(ready_o),
        .data_i(data_i),
        .data_a_o(ram_row0),
        .data_b_o(ram_row1)
    );

    // convolution sliding window
    logic [WIDTH_P-1:0] conv_window [2:0][2:0];

    integer r;
    integer c;

    always_ff @(posedge clk_i) begin
        if (!rstn_i) begin
            for (r = 0; r < 3; r = r + 1) begin
                for (c = 0; c < 3; c = c + 1) begin
                    conv_window[r][c] <= '0;
                end
            end
        end else if (valid_i & ready_o) begin
            // shift data into each row
            for (r = 0; r < 3; r = r + 1) begin
                conv_window[r][0] <= conv_window[r][1];
                conv_window[r][1] <= conv_window[r][2];
            end
            
            // shift corresponding row data into each row
            conv_window[0][2] <= ram_row0; // 2 rows ago
            conv_window[1][2] <= ram_row1; // 1 row ago
            conv_window[2][2] <= data_i; // newest data
        end
    end

    // sobel x and y kernel
    // 1d 2d arrays not supported in icarus???
    // localparam signed [3:0] KX [8:0] = '{
    //     -1,  0,  1,
    //     -2,  0,  2,
    //     -1,  0,  1
    // };
    
    // localparam signed [3:0] KY [8:0] = '{
    //     -1, -2, -1,
    //      0,  0,  0,
    //      1,  2,  1
    // };
    function automatic signed [3:0] kx;
        input integer idx;
        begin
            case (idx)
                0: kx = -1;  1: kx =  0;  2: kx =  1;
                3: kx = -2;  4: kx =  0;  5: kx =  2;
                6: kx = -1;  7: kx =  0;  8: kx =  1;
                default: kx = 0;
            endcase
        end
    endfunction

    function automatic signed [3:0] ky;
        input integer idx;
        begin
            case (idx)
                0: ky = -1;  1: ky = -2;  2: ky = -1;
                3: ky =  0;  4: ky =  0;  5: ky =  0;
                6: ky =  1;  7: ky =  2;  8: ky =  1;
                default: ky = 0;
            endcase
        end
    endfunction

    logic signed [(2*WIDTH_P)-1:0] gx_sum [0:8];
    logic signed [(2*WIDTH_P)-1:0] gy_sum [0:8];

    assign gx_sum[0] = $signed({1'b0, conv_window[0][0]}) * kx(0);
    assign gy_sum[0] = $signed({1'b0, conv_window[0][0]}) * ky(0);

    genvar t;
    generate
        for (t = 1; t < 9; t = t + 1) begin
            // converted to unsigned to match the jupyter model
            assign gx_sum[t] = gx_sum[t-1] + ($signed({1'b0, conv_window[t/3][t%3]}) * kx(t)); // v*erilator wants to flatten this so it gives a circular comb error but its an prefix counter so its expected
            assign gy_sum[t] = gy_sum[t-1] + ($signed({1'b0, conv_window[t/3][t%3]}) * ky(t));
        end
    endgenerate

    // gradient is sum of all previous values
    assign gx_o = gx_sum[8];
    assign gy_o = gy_sum[8];
endmodule
