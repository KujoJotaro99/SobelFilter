`timescale 1ns/1ps

module rgb2gray_tb;
endmodule
