`timescale 1ns/1ps

module sobel (
);
endmodule
