module spi_axis (
);
endmodule
